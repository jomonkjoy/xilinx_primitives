
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
//     19-36      |  "36Kb"   |    1024   |    10-bit     |    4-bit    //
//     10-18      |  "36Kb"   |    2048   |    11-bit     |    2-bit    //
//     10-18      |  "18Kb"   |    1024   |    10-bit     |    2-bit    //
//      5-9       |  "36Kb"   |    4096   |    12-bit     |    1-bit    //
//      5-9       |  "18Kb"   |    2048   |    11-bit     |    1-bit    //
//      3-4       |  "36Kb"   |    8192   |    13-bit     |    1-bit    //
//      3-4       |  "18Kb"   |    4096   |    12-bit     |    1-bit    //
//        2       |  "36Kb"   |   16384   |    14-bit     |    1-bit    //
//        2       |  "18Kb"   |    8192   |    13-bit     |    1-bit    //
//        1       |  "36Kb"   |   32768   |    15-bit     |    1-bit    //
//        1       |  "18Kb"   |   16384   |    14-bit     |    1-bit    //
//////////////////////////////////////////////////////////////////////////

module xilinx_tdp_bram 
import xilinx_primitive_pkg::*;
#(
   parameter BRAM_SIZE              = "18Kb", // Target BRAM: "18Kb" or "36Kb"
   parameter DEVICE                 = "7SERIES", // Target device: "7SERIES"
   parameter DOA_REG                = 0,        // Optional port A output register (0 or 1)
   parameter DOB_REG                = 0,        // Optional port B output register (0 or 1)
   parameter INIT_A                 = 36'h0000000,  // Initial values on port A output port
   parameter INIT_B                 = 36'h00000000, // Initial values on port B output port
   parameter INIT_FILE              = "NONE",
   parameter READ_WIDTH_A           = 1,   // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
   parameter READ_WIDTH_B           = 1,   // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
   parameter SIM_COLLISION_CHECK    = "ALL", // Collision check enable "ALL", "WARNING_ONLY",
                                            //   "GENERATE_X_ONLY" or "NONE"
   parameter SRVAL_A                = 36'h00000000, // Set/Reset value for port A output
   parameter SRVAL_B                = 36'h00000000, // Set/Reset value for port B output
   parameter WRITE_MODE_A           = "WRITE_FIRST", // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
   parameter WRITE_MODE_B           = "WRITE_FIRST", // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
   parameter WRITE_WIDTH_A          = 1, // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
   parameter WRITE_WIDTH_B          = 1  // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
) (
   output logic [READ_WIDTH_A-1:0]  DOA,       // Output port-A data, width defined by READ_WIDTH_A parameter
   output logic [READ_WIDTH_B-1:0]  DOB,       // Output port-B data, width defined by READ_WIDTH_B parameter
   input  logic [14:0]              ADDRA,     // Input port-A address, width defined by Port A depth
   input  logic [14:0]              ADDRB,     // Input port-B address, width defined by Port B depth
   input  logic                     CLKA,      // 1-bit input port-A clock
   input  logic                     CLKB,      // 1-bit input port-B clock
   input  logic [WRITE_WIDTH_A-1:0] DIA,       // Input port-A data, width defined by WRITE_WIDTH_A parameter
   input  logic [WRITE_WIDTH_B-1:0] DIB,       // Input port-B data, width defined by WRITE_WIDTH_B parameter
   input  logic                     ENA,       // 1-bit input port-A enable
   input  logic                     ENB,       // 1-bit input port-B enable
   input  logic                     REGCEA,    // 1-bit input port-A output register enable
   input  logic                     REGCEB,    // 1-bit input port-B output register enable
   input  logic                     RSTA,      // 1-bit input port-A reset
   input  logic                     RSTB,      // 1-bit input port-B reset
   input  logic [3:0]               WEA,       // Input port-A write enable, width defined by Port A depth
   input  logic [3:0]               WEB        // Input port-B write enable, width defined by Port B depth
);

localparam MACRO_SIZE = (WRITE_WIDTH_A>16 || WRITE_WIDTH_B>16) ? "36Kb" : BRAM_SIZE;
localparam BRAM_DEPTH_A = get_tdp_bram_depth(WRITE_WIDTH_A, MACRO_SIZE);
localparam BRAM_DEPTH_B = get_tdp_bram_depth(WRITE_WIDTH_B, MACRO_SIZE);
localparam BRAM_WE_A = get_tdp_we_width(WRITE_WIDTH_A);
localparam BRAM_WE_B = get_tdp_we_width(WRITE_WIDTH_B);
localparam ADDR_WIDTH_A = $clog2(BRAM_DEPTH_A);
localparam ADDR_WIDTH_B = $clog2(BRAM_DEPTH_B);

generate if (MACRO_SIZE=="18Kb") begin

// Internal signals for RAMB18E1
logic [15:0] DOADO_wire;
logic [15:0] DOBDO_wire;
logic [1:0]  DOPADOP_wire;
logic [1:0]  DOPBDOP_wire;
logic [13:0] ADDRARDADDR_wire;
logic [13:0] ADDRBWRADDR_wire;
logic [15:0] DIADI_wire;
logic [15:0] DIBDI_wire;
logic [1:0]  DIPADIP_wire;
logic [1:0]  DIPBDIP_wire;
logic [1:0]  WEA_wire;
logic [3:0]  WEBWE_wire;

// Address mapping for 18Kb BRAM (14-bit address bus)
assign ADDRARDADDR_wire = {{(14-ADDR_WIDTH_A){1'b0}}, ADDRA[ADDR_WIDTH_A-1:0]};
assign ADDRBWRADDR_wire = {{(14-ADDR_WIDTH_B){1'b0}}, ADDRB[ADDR_WIDTH_B-1:0]};
   
// Data input mapping
assign DIADI_wire = {{(16-WRITE_WIDTH_A){1'b0}}, DIA};
assign DIBDI_wire = {{(16-WRITE_WIDTH_B){1'b0}}, DIB};
assign DIPADIP_wire = 2'b00;
assign DIPBDIP_wire = 2'b00;
   
// Data output mapping
assign DOA = DOADO_wire[READ_WIDTH_A-1:0];
assign DOB = DOBDO_wire[READ_WIDTH_B-1:0];
   
// Write enable mapping
assign WEA_wire = WEA[BRAM_WE_A-1:0];
assign WEBWE_wire = {2'b00, WEB[BRAM_WE_B-1:0]};

// RAMB18E1: 18K-bit Configurable Synchronous Block RAM
//           7 Series
// Xilinx HDL Language Template, version 2025.1

RAMB18E1 #(
   // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
   .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
   // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
   .SIM_COLLISION_CHECK("ALL"),
   // DOA_REG, DOB_REG: Optional output register (0 or 1)
   .DOA_REG(DOA_REG),
   .DOB_REG(DOB_REG),
   // INITP_00 to INITP_07: Initial contents of parity memory array
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_00 to INIT_3F: Initial contents of data memory array
   .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_A, INIT_B: Initial values on output ports
   .INIT_A(18'h00000),
   .INIT_B(18'h00000),
   // Initialization File: RAM initialization file
   .INIT_FILE("NONE"),
   // RAM Mode: "SDP" or "TDP"
   .RAM_MODE("TDP"),
   // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
   .READ_WIDTH_A(READ_WIDTH_A),                                                                 // 0-72
   .READ_WIDTH_B(READ_WIDTH_B),                                                                 // 0-18
   .WRITE_WIDTH_A(WRITE_WIDTH_A),                                                               // 0-18
   .WRITE_WIDTH_B(WRITE_WIDTH_B),                                                               // 0-72
   // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
   .RSTREG_PRIORITY_A("RSTREG"),
   .RSTREG_PRIORITY_B("RSTREG"),
   // SRVAL_A, SRVAL_B: Set/reset value for output
   .SRVAL_A(18'h00000),
   .SRVAL_B(18'h00000),
   // Simulation Device: Must be set to "7SERIES" for simulation behavior
   .SIM_DEVICE("7SERIES"),
   // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
   .WRITE_MODE_A(WRITE_MODE_A),
   .WRITE_MODE_B(WRITE_MODE_B)
)
RAMB18E1_inst (
   // Port A Data: 16-bit (each) output: Port A data
   .DOADO(DOADO_wire),            // 16-bit output: A port data/LSB data
   .DOPADOP(DOPADOP_wire),        // 2-bit output: A port parity/LSB parity
   // Port B Data: 16-bit (each) output: Port B data
   .DOBDO(DOBDO_wire),            // 16-bit output: B port data/MSB data
   .DOPBDOP(DOPBDOP_wire),        // 2-bit output: B port parity/MSB parity
   // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
   // when RAM_MODE="SDP")
   .ADDRARDADDR(ADDRARDADDR_wire),// 14-bit input: A port address/Read address
   .CLKARDCLK(CLKA),              // 1-bit input: A port clock/Read clock
   .ENARDEN(ENA),                 // 1-bit input: A port enable/Read enable
   .REGCEAREGCE(REGCEA),          // 1-bit input: A port register enable/Register enable
   .RSTRAMARSTRAM(RSTA),          // 1-bit input: A port set/reset
   .RSTREGARSTREG(RSTA),          // 1-bit input: A port register set/reset
   .WEA(WEA_wire),                // 2-bit input: A port write enable
   // Port A Data: 16-bit (each) input: Port A data
   .DIADI(DIADI_wire),            // 16-bit input: A port data/LSB data
   .DIPADIP(DIPADIP_wire),        // 2-bit input: A port parity/LSB parity
   // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
   // when RAM_MODE="SDP")
   .ADDRBWRADDR(ADDRBWRADDR_wire),// 14-bit input: B port address/Write address
   .CLKBWRCLK(CLKB),              // 1-bit input: B port clock/Write clock
   .ENBWREN(ENB),                 // 1-bit input: B port enable/Write enable
   .REGCEB(REGCEB),               // 1-bit input: B port register enable
   .RSTRAMB(RSTB),                // 1-bit input: B port set/reset
   .RSTREGB(RSTB),                // 1-bit input: B port register set/reset
   .WEBWE(WEBWE_wire),            // 4-bit input: B port write enable/Write enable
   // Port B Data: 16-bit (each) input: Port B data
   .DIBDI(DIBDI_wire),            // 16-bit input: B port data/MSB data
   .DIPBDIP(DIPBDIP_wire)         // 2-bit input: B port parity/MSB parity
);

// End of RAMB18E1_inst instantiation

end else begin

// Internal signals for RAMB36E1
logic [31:0] DOADO_wire;
logic [31:0] DOBDO_wire;
logic [3:0]  DOPADOP_wire;
logic [3:0]  DOPBDOP_wire;
logic [15:0] ADDRARDADDR_wire;
logic [15:0] ADDRBWRADDR_wire;
logic [31:0] DIADI_wire;
logic [31:0] DIBDI_wire;
logic [3:0]  DIPADIP_wire;
logic [3:0]  DIPBDIP_wire;
logic [3:0]  WEA_wire;
logic [7:0]  WEBWE_wire;

// Address mapping for 36Kb BRAM (16-bit address bus)
assign ADDRARDADDR_wire = {{(16-ADDR_WIDTH_A){1'b0}}, ADDRA[ADDR_WIDTH_A-1:0]};
assign ADDRBWRADDR_wire = {{(16-ADDR_WIDTH_B){1'b0}}, ADDRB[ADDR_WIDTH_B-1:0]};
   
// Data input mapping
assign DIADI_wire = {{(32-WRITE_WIDTH_A){1'b0}}, DIA};
assign DIBDI_wire = {{(32-WRITE_WIDTH_B){1'b0}}, DIB};
assign DIPADIP_wire = 4'b0000;
assign DIPBDIP_wire = 4'b0000;
   
// Data output mapping
assign DOA = DOADO_wire[READ_WIDTH_A-1:0];
assign DOB = DOBDO_wire[READ_WIDTH_B-1:0];
   
// Write enable mapping
assign WEA_wire = {{(4-BRAM_WE_A){1'b0}}, WEA[BRAM_WE_A-1:0]};
assign WEBWE_wire = {{(4-BRAM_WE_B){1'b0}}, WEB[BRAM_WE_B-1:0], 4'b0000};

// RAMB36E1: 36K-bit Configurable Synchronous Block RAM
//           7 Series
// Xilinx HDL Language Template, version 2025.1

RAMB36E1 #(
   // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
   .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
   // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
   .SIM_COLLISION_CHECK("ALL"),
   // DOA_REG, DOB_REG: Optional output register (0 or 1)
   .DOA_REG(DOA_REG),
   .DOB_REG(DOB_REG),
   .EN_ECC_READ("FALSE"),                                                            // Enable ECC decoder,
                                                                                     // FALSE, TRUE
   .EN_ECC_WRITE("FALSE"),                                                           // Enable ECC encoder,
                                                                                     // FALSE, TRUE
   // INITP_00 to INITP_0F: Initial contents of the parity memory array
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_00 to INIT_7F: Initial contents of the data memory array
   .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_A, INIT_B: Initial values on output ports
   .INIT_A(36'h000000000),
   .INIT_B(36'h000000000),
   // Initialization File: RAM initialization file
   .INIT_FILE("NONE"),
   // RAM Mode: "SDP" or "TDP"
   .RAM_MODE("TDP"),
   // RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
   .RAM_EXTENSION_A("NONE"),
   .RAM_EXTENSION_B("NONE"),
   // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
   .READ_WIDTH_A(READ_WIDTH_A),                                                                 // 0-72
   .READ_WIDTH_B(READ_WIDTH_B),                                                                 // 0-36
   .WRITE_WIDTH_A(WRITE_WIDTH_A),                                                               // 0-36
   .WRITE_WIDTH_B(WRITE_WIDTH_B),                                                               // 0-72
   // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
   .RSTREG_PRIORITY_A("RSTREG"),
   .RSTREG_PRIORITY_B("RSTREG"),
   // SRVAL_A, SRVAL_B: Set/reset value for output
   .SRVAL_A(36'h000000000),
   .SRVAL_B(36'h000000000),
   // Simulation Device: Must be set to "7SERIES" for simulation behavior
   .SIM_DEVICE("7SERIES"),
   // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
   .WRITE_MODE_A(WRITE_MODE_A),
   .WRITE_MODE_B(WRITE_MODE_B)
)
RAMB36E1_inst (
   // Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
   .CASCADEOUTA(),                // 1-bit output: A port cascade
   .CASCADEOUTB(),                // 1-bit output: B port cascade
   // ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
   .DBITERR(),                    // 1-bit output: Double bit error status
   .ECCPARITY(),                  // 8-bit output: Generated error correction parity
   .RDADDRECC(),                  // 9-bit output: ECC read address
   .SBITERR(),                    // 1-bit output: Single bit error status
   // Port A Data: 32-bit (each) output: Port A data
   .DOADO(DOADO_wire),            // 32-bit output: A port data/LSB data
   .DOPADOP(DOPADOP_wire),        // 4-bit output: A port parity/LSB parity
   // Port B Data: 32-bit (each) output: Port B data
   .DOBDO(DOBDO_wire),            // 32-bit output: B port data/MSB data
   .DOPBDOP(DOPBDOP_wire),        // 4-bit output: B port parity/MSB parity
   // Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
   .CASCADEINA(0),                // 1-bit input: A port cascade
   .CASCADEINB(0),                // 1-bit input: B port cascade
   // ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
   .INJECTDBITERR(0),             // 1-bit input: Inject a double bit error
   .INJECTSBITERR(0),             // 1-bit input: Inject a single bit error
   // Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
   // when RAM_MODE="SDP")
   .ADDRARDADDR(ADDRARDADDR_wire),// 16-bit input: A port address/Read address
   .CLKARDCLK(CLKA),              // 1-bit input: A port clock/Read clock
   .ENARDEN(ENA),                 // 1-bit input: A port enable/Read enable
   .REGCEAREGCE(REGCEA),          // 1-bit input: A port register enable/Register enable
   .RSTRAMARSTRAM(RSTA),          // 1-bit input: A port set/reset
   .RSTREGARSTREG(RSTA),          // 1-bit input: A port register set/reset
   .WEA(WEA_wire),                // 4-bit input: A port write enable
   // Port A Data: 32-bit (each) input: Port A data
   .DIADI(DIADI_wire),            // 32-bit input: A port data/LSB data
   .DIPADIP(DIPADIP_wire),        // 4-bit input: A port parity/LSB parity
   // Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
   // when RAM_MODE="SDP")
   .ADDRBWRADDR(ADDRBWRADDR_wire),// 16-bit input: B port address/Write address
   .CLKBWRCLK(CLKB),              // 1-bit input: B port clock/Write clock
   .ENBWREN(ENB),                 // 1-bit input: B port enable/Write enable
   .REGCEB(REGCEB),               // 1-bit input: B port register enable
   .RSTRAMB(RSTB),                // 1-bit input: B port set/reset
   .RSTREGB(RSTB),                // 1-bit input: B port register set/reset
   .WEBWE(WEBWE_wire),            // 8-bit input: B port write enable/Write enable
   // Port B Data: 32-bit (each) input: Port B data
   .DIBDI(DIBDI_wire),            // 32-bit input: B port data/MSB data
   .DIPBDIP(DIPBDIP_wire)         // 4-bit input: B port parity/MSB parity
);

// End of RAMB36E1_inst instantiation

end endgenerate

endmodule
