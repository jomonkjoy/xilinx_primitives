
///////////////////////////////////////////////////////////////////////
//  READ_WIDTH | BRAM_SIZE | READ Depth  | RDADDR Width |            //
// WRITE_WIDTH |           | WRITE Depth | WRADDR Width |  WE Width  //
// ============|===========|=============|==============|============//
//    37-72    |  "36Kb"   |      512    |     9-bit    |    8-bit   //
//    19-36    |  "36Kb"   |     1024    |    10-bit    |    4-bit   //
//    19-36    |  "18Kb"   |      512    |     9-bit    |    4-bit   //
//    10-18    |  "36Kb"   |     2048    |    11-bit    |    2-bit   //
//    10-18    |  "18Kb"   |     1024    |    10-bit    |    2-bit   //
//     5-9     |  "36Kb"   |     4096    |    12-bit    |    1-bit   //
//     5-9     |  "18Kb"   |     2048    |    11-bit    |    1-bit   //
//     3-4     |  "36Kb"   |     8192    |    13-bit    |    1-bit   //
//     3-4     |  "18Kb"   |     4096    |    12-bit    |    1-bit   //
//       2     |  "36Kb"   |    16384    |    14-bit    |    1-bit   //
//       2     |  "18Kb"   |     8192    |    13-bit    |    1-bit   //
//       1     |  "36Kb"   |    32768    |    15-bit    |    1-bit   //
//       1     |  "18Kb"   |    16384    |    14-bit    |    1-bit   //
///////////////////////////////////////////////////////////////////////

module xilinx_sdp_bram 
import xilinx_primitive_pkg::*;
#(
   parameter BRAM_SIZE              = "18Kb", // Target BRAM, "18Kb" or "36Kb"
   parameter DEVICE                 = "7SERIES", // Target device: "7SERIES"
   parameter WRITE_WIDTH            = 1,        // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
   parameter READ_WIDTH             = 1,        // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
   parameter DO_REG                 = 0,        // Optional output register (0 or 1)
   parameter INIT_FILE              = "NONE",
   parameter SIM_COLLISION_CHECK    = "ALL",    // Collision check enable "ALL", "WARNING_ONLY",
                                                //   "GENERATE_X_ONLY" or "NONE"
   parameter SRVAL                  = 72'h000000000000000000, // Set/Reset value for port output
   parameter INIT                   = 72'h000000000000000000,  // Initial values on output port
   parameter WRITE_MODE             = "WRITE_FIRST"  // Specify "READ_FIRST" for same clock or synchronous clocks
                                                    //   Specify "WRITE_FIRST for asynchronous clocks on ports
) (
   output logic [READ_WIDTH-1:0]    DO,         // Output read data port, width defined by READ_WIDTH parameter
   input  logic [WRITE_WIDTH-1:0]   DI,         // Input write data port, width defined by WRITE_WIDTH parameter
   input  logic [14:0]              RDADDR,     // Input read address, width defined by read port depth
   input  logic                     RDCLK,      // 1-bit input read clock
   input  logic                     RDEN,       // 1-bit input read port enable
   input  logic                     REGCE,      // 1-bit input read output register enable
   input  logic                     RST,        // 1-bit input reset
   input  logic [7:0]               WE,         // Input write enable, width defined by write port depth
   input  logic [14:0]              WRADDR,     // Input write address, width defined by write port depth
   input  logic                     WRCLK,      // 1-bit input write clock
   input  logic                     WREN        // 1-bit input write port enable
);

localparam MACRO_SIZE = (WRITE_WIDTH>32) ? "36Kb" : BRAM_SIZE;
localparam WRITE_DEPTH = get_sdp_depth(WRITE_WIDTH, BRAM_SIZE);
localparam READ_DEPTH = get_sdp_depth(READ_WIDTH, BRAM_SIZE);
localparam BRAM_WE = get_sdp_we_width(WRITE_WIDTH);

// Calculate address widths based on depth
localparam WRADDR_WIDTH = $clog2(WRITE_DEPTH);
localparam RDADDR_WIDTH = $clog2(READ_DEPTH);

// Internal signals for BRAM primitives
logic [31:0] DOADO_wire;
logic [3:0]  DOPADOP_wire;
logic [31:0] DIBDI_wire;
logic [3:0]  DIPBDIP_wire;
logic [15:0] ADDRARDADDR_wire;
logic [15:0] ADDRBWRADDR_wire;
logic [7:0]  WEBWE_wire;

// Address adjustment - BRAM addresses are word-aligned
// For 18Kb BRAM: ADDR[13:0], for 36Kb BRAM: ADDR[15:0]
always_comb begin
   // Read address - adjust based on data width
   if (READ_WIDTH <= 1)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:0]};
   else if (READ_WIDTH <= 2)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:1], 1'b0};
   else if (READ_WIDTH <= 4)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:2], 2'b00};
   else if (READ_WIDTH <= 9)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:3], 3'b000};
   else if (READ_WIDTH <= 18)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:4], 4'b0000};
   else if (READ_WIDTH <= 36)
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:5], 5'b00000};
   else // 37-72
      ADDRARDADDR_wire = {1'b1, RDADDR[RDADDR_WIDTH-1:6], 6'b000000};
      
   // Write address - adjust based on data width
   if (WRITE_WIDTH <= 1)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:0]};
   else if (WRITE_WIDTH <= 2)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:1], 1'b0};
   else if (WRITE_WIDTH <= 4)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:2], 2'b00};
   else if (WRITE_WIDTH <= 9)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:3], 3'b000};
   else if (WRITE_WIDTH <= 18)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:4], 4'b0000};
   else if (WRITE_WIDTH <= 36)
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:5], 5'b00000};
   else // 37-72
      ADDRBWRADDR_wire = {1'b1, WRADDR[WRADDR_WIDTH-1:6], 6'b000000};
end

// Data input mapping
assign DIBDI_wire = {{(32-WRITE_WIDTH){1'b0}}, DI};
assign DIPBDIP_wire = 4'b0000;
   
// Data output mapping
assign DO = DOADO_wire[READ_WIDTH-1:0];
   
// Write enable mapping
assign WEBWE_wire = {{(4-BRAM_WE){1'b0}}, WE[BRAM_WE-1:0]};

generate if (MACRO_SIZE=="18Kb") begin

// RAMB18E1: 18K-bit Configurable Synchronous Block RAM
//           7 Series
// Xilinx HDL Language Template, version 2025.1

RAMB18E1 #(
   // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
   .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
   // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
   .SIM_COLLISION_CHECK("ALL"),
   // DOA_REG, DOB_REG: Optional output register (0 or 1)
   .DOA_REG(0),
   .DOB_REG(0),
   // INITP_00 to INITP_07: Initial contents of parity memory array
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_00 to INIT_3F: Initial contents of data memory array
   .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_A, INIT_B: Initial values on output ports
   .INIT_A(18'h00000),
   .INIT_B(18'h00000),
   // Initialization File: RAM initialization file
   .INIT_FILE("NONE"),
   // RAM Mode: "SDP" or "TDP"
   .RAM_MODE("SDP"),
   // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
   .READ_WIDTH_A(READ_WIDTH),                                                        // 0-72
   .READ_WIDTH_B(0),                                                                 // 0-18
   .WRITE_WIDTH_A(0),                                                                // 0-18
   .WRITE_WIDTH_B(WRITE_WIDTH),                                                      // 0-72
   // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
   .RSTREG_PRIORITY_A("RSTREG"),
   .RSTREG_PRIORITY_B("RSTREG"),
   // SRVAL_A, SRVAL_B: Set/reset value for output
   .SRVAL_A(18'h00000),
   .SRVAL_B(18'h00000),
   // Simulation Device: Must be set to "7SERIES" for simulation behavior
   .SIM_DEVICE("7SERIES"),
   // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
   .WRITE_MODE_A("NO_CHANGE"),
   .WRITE_MODE_B(WRITE_MODE)
)
RAMB18E1_inst (
   // Port A Data: 16-bit (each) output: Port A data
   .DOADO(DOADO_wire[15:0]),      // 16-bit output: A port data/LSB data
   .DOPADOP(DOPADOP_wire[1:0]),   // 2-bit output: A port parity/LSB parity
   // Port B Data: 16-bit (each) output: Port B data
   .DOBDO(),                      // 16-bit output: B port data/MSB data
   .DOPBDOP(),                    // 2-bit output: B port parity/MSB parity
   // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
   // when RAM_MODE="SDP")
   .ADDRARDADDR(ADDRARDADDR_wire[13:0]),// 14-bit input: A port address/Read address
   .CLKARDCLK(RDCLK),             // 1-bit input: A port clock/Read clock
   .ENARDEN(RDEN),                // 1-bit input: A port enable/Read enable
   .REGCEAREGCE(REGCE),           // 1-bit input: A port register enable/Register enable
   .RSTRAMARSTRAM(RST),           // 1-bit input: A port set/reset
   .RSTREGARSTREG(RST),           // 1-bit input: A port register set/reset
   .WEA(0),                       // 2-bit input: A port write enable
   // Port A Data: 16-bit (each) input: Port A data
   .DIADI(0),                     // 16-bit input: A port data/LSB data
   .DIPADIP(0),                   // 2-bit input: A port parity/LSB parity
   // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
   // when RAM_MODE="SDP")
   .ADDRBWRADDR(ADDRBWRADDR_wire[13:0]),// 14-bit input: B port address/Write address
   .CLKBWRCLK(WRCLK),             // 1-bit input: B port clock/Write clock
   .ENBWREN(WREN),                // 1-bit input: B port enable/Write enable
   .REGCEB(0),                    // 1-bit input: B port register enable
   .RSTRAMB(RST),                 // 1-bit input: B port set/reset
   .RSTREGB(RST),                 // 1-bit input: B port register set/reset
   .WEBWE(WEBWE_wire[3:0]),       // 4-bit input: B port write enable/Write enable
   // Port B Data: 16-bit (each) input: Port B data
   .DIBDI(DIBDI_wire[15:0]),      // 16-bit input: B port data/MSB data
   .DIPBDIP(DIPBDIP_wire[1:0])    // 2-bit input: B port parity/MSB parity
);

// End of RAMB18E1_inst instantiation

end else begin

// RAMB36E1: 36K-bit Configurable Synchronous Block RAM
//           7 Series
// Xilinx HDL Language Template, version 2025.1

RAMB36E1 #(
   // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
   .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
   // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
   .SIM_COLLISION_CHECK("ALL"),
   // DOA_REG, DOB_REG: Optional output register (0 or 1)
   .DOA_REG(0),
   .DOB_REG(0),
   .EN_ECC_READ("FALSE"),                                                            // Enable ECC decoder,
                                                                                     // FALSE, TRUE
   .EN_ECC_WRITE("FALSE"),                                                           // Enable ECC encoder,
                                                                                     // FALSE, TRUE
   // INITP_00 to INITP_0F: Initial contents of the parity memory array
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_00 to INIT_7F: Initial contents of the data memory array
   .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_A, INIT_B: Initial values on output ports
   .INIT_A(36'h000000000),
   .INIT_B(36'h000000000),
   // Initialization File: RAM initialization file
   .INIT_FILE("NONE"),
   // RAM Mode: "SDP" or "TDP"
   .RAM_MODE("SDP"),
   // RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
   .RAM_EXTENSION_A("NONE"),
   .RAM_EXTENSION_B("NONE"),
   // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
   .READ_WIDTH_A(READ_WIDTH),                                                        // 0-72
   .READ_WIDTH_B(0),                                                                 // 0-36
   .WRITE_WIDTH_A(0),                                                                // 0-36
   .WRITE_WIDTH_B(WRITE_WIDTH),                                                      // 0-72
   // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
   .RSTREG_PRIORITY_A("RSTREG"),
   .RSTREG_PRIORITY_B("RSTREG"),
   // SRVAL_A, SRVAL_B: Set/reset value for output
   .SRVAL_A(36'h000000000),
   .SRVAL_B(36'h000000000),
   // Simulation Device: Must be set to "7SERIES" for simulation behavior
   .SIM_DEVICE("7SERIES"),
   // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
   .WRITE_MODE_A("NO_CHANGE"),
   .WRITE_MODE_B(WRITE_MODE)
)
RAMB36E1_inst (
   // Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
   .CASCADEOUTA(),                // 1-bit output: A port cascade
   .CASCADEOUTB(),                // 1-bit output: B port cascade
   // ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
   .DBITERR(),                    // 1-bit output: Double bit error status
   .ECCPARITY(),                  // 8-bit output: Generated error correction parity
   .RDADDRECC(),                  // 9-bit output: ECC read address
   .SBITERR(),                    // 1-bit output: Single bit error status
   // Port A Data: 32-bit (each) output: Port A data
   .DOADO(DOADO_wire[31:0]),      // 32-bit output: A port data/LSB data
   .DOPADOP(DOPADOP_wire[3:0]),   // 4-bit output: A port parity/LSB parity
   // Port B Data: 32-bit (each) output: Port B data
   .DOBDO(),                      // 32-bit output: B port data/MSB data
   .DOPBDOP(),                    // 4-bit output: B port parity/MSB parity
   // Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
   .CASCADEINA(0),                // 1-bit input: A port cascade
   .CASCADEINB(0),                // 1-bit input: B port cascade
   // ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
   .INJECTDBITERR(0),             // 1-bit input: Inject a double bit error
   .INJECTSBITERR(0),             // 1-bit input: Inject a single bit error
   // Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
   // when RAM_MODE="SDP")
   .ADDRARDADDR(ADDRARDADDR_wire[15:0]),// 16-bit input: A port address/Read address
   .CLKARDCLK(RDCLK),             // 1-bit input: A port clock/Read clock
   .ENARDEN(RDEN),                // 1-bit input: A port enable/Read enable
   .REGCEAREGCE(REGCE),           // 1-bit input: A port register enable/Register enable
   .RSTRAMARSTRAM(RST),           // 1-bit input: A port set/reset
   .RSTREGARSTREG(RST),           // 1-bit input: A port register set/reset
   .WEA(0),                       // 4-bit input: A port write enable
   // Port A Data: 32-bit (each) input: Port A data
   .DIADI(0),                     // 32-bit input: A port data/LSB data
   .DIPADIP(0),                   // 4-bit input: A port parity/LSB parity
   // Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
   // when RAM_MODE="SDP")
   .ADDRBWRADDR(ADDRBWRADDR_wire[15:0]),// 16-bit input: B port address/Write address
   .CLKBWRCLK(WRCLK),             // 1-bit input: B port clock/Write clock
   .ENBWREN(WREN),                // 1-bit input: B port enable/Write enable
   .REGCEB(0),                    // 1-bit input: B port register enable
   .RSTRAMB(RST),                 // 1-bit input: B port set/reset
   .RSTREGB(RST),                 // 1-bit input: B port register set/reset
   .WEBWE(WEBWE_wire[7:0]),       // 8-bit input: B port write enable/Write enable
   // Port B Data: 32-bit (each) input: Port B data
   .DIBDI(DIBDI_wire[31:0]),      // 32-bit input: B port data/MSB data
   .DIPBDIP(DIPBDIP_wire[3:0])    // 4-bit input: B port parity/MSB parity
);

// End of RAMB36E1_inst instantiation

end endgenerate

endmodule
